magic
tech scmos
timestamp 1763640429
<< nwell >>
rect -1 6 30 18
<< polysilicon >>
rect 7 17 10 19
rect 18 17 21 19
rect 7 2 10 7
rect -1 -1 10 2
rect 7 -6 10 -1
rect 18 5 21 7
rect 18 2 31 5
rect 18 -6 21 2
rect 7 -19 10 -17
rect 18 -19 21 -17
<< ndiffusion >>
rect 0 -17 7 -6
rect 10 -17 18 -6
rect 21 -17 31 -6
<< pdiffusion >>
rect 0 7 7 17
rect 10 7 18 17
rect 21 7 29 17
<< metal1 >>
rect -2 24 31 29
rect 1 8 6 24
rect 12 0 17 16
rect 23 8 28 24
rect 12 -3 39 0
rect 1 -23 6 -8
rect 24 -15 29 -3
rect 1 -27 31 -23
<< ntransistor >>
rect 7 -17 10 -6
rect 18 -17 21 -6
<< ptransistor >>
rect 7 7 10 17
rect 18 7 21 17
<< labels >>
rlabel polysilicon 0 -1 8 1 1 a
rlabel polysilicon 23 3 31 5 1 b
rlabel metal1 14 -26 22 -24 1 gnd
rlabel metal1 13 26 21 28 5 vdd
rlabel metal1 31 -2 39 0 7 out
<< end >>
